OEMs/BPTvJyz56VSjS4kxHdkYM07ab9x+
e5lfzcLobINV4xvCgWeB1d4Z13gakeqSnX3fP342f73QTa8eGkfaNSzgCiH7gT5FDI+cBZCfPnFU
a4NoorrIulQ2fZKgMIN95eD/jJ3p2nI1QDaPOiSDNvsnnrk50YXTapUvQODp90zMTRg0ZUHalNwg
TiDGzR/oVpwNxUAQgEsLeVHrff8p8UKSRWI6RJ926Ogl5LV2HDNCQYwWEpGokaboQRAY310PSWI6
pBMcwZipLoFwkBIynZW7ZvKYt4aGZUf5vgfAB1MxftQ1hNvJ+sgEPBSAH2ibSGPjdkI2bXvRRCvv
RG7o6LoEiSW9M/7xXTz7T6l+QrIIyu+YZiKwX7/xQGBN8Clx5GFJI8QF/wPNeFwnjD98ZvNxL4tK
/PYBEt03+IkxL9Aozvj6DDKZNvetDcBIksKQ/fIpqUEisRX7C/4paddKwwMaf+yMICcAqcTCSChM
TrjWROqPl4afwyZHMEUfQlu0fGxB+bqN+uzVVQdq8uz9s+nlFkkm/eKgX+1YjTCewiO4wWMPC4KF
dj6vxxcig4jIx5b6wM3tcFxpavIY+Q2VWQwg8ZFR0pf3x3vcAQclSlGBDAgvknJGisEbKLIYq+SL
HoxtlyGtuhRRjCsGngabAfceqiNiG1Bxu8sIqVmlrQQjWBXMAG1zoEUMvyAFpMtFgTiaabjPEjvZ
9/KUM2GeTRVNbcxJzaeU09HPkV/u/KghqtfLtzF+dvct+G6lrh1iISXKXu8E8NpYNjkcKMuasbdU
Yy4Ew7z3C7YC1Y8Gm8/inWvolc/Zgf+n9U8GlzxtnIXF5lJHbUKrKjOW06krHNp/kOjiZcQ/HZ5F
npYzFPSl7+7FcaQVWuUYpHBWJwA737AY3Pd9GrvciGgjnCIe4Dt+DWRWQM5PbReJjdpFq5d9RSbK
oycW4XyJwzu3J4HDhJLT9hwD6mVt9uOWp6P0qn5vginxtfaYOQwlIL7OrjwE0xto1xtNAP+ngQJm
jTwwbb/TDuE5Cokd4IWGA9vMyWO5l1J1SkWM55mu8W+2VDsUA9pQ0gcs6K+PlBw0d0QO2ejF8o9r
vj7ggmSAHKAA+/T3RGJIFKBFscxRR11+VZj9VUL9TNKTg/A2p/qCPwDA3azuYoCH7vhAUi2Z+zzQ
WuS+YsU2XtkGeTY7FMd58b1/lUXwL6S5R6ej8ZkSVztU25rtaKWZFotQnP65zFGlx9oVqdha8MgU
rnlWDc106gDzJ/C27uX+B2vby/jlS1KFpJ1BhFoTRmoOscFWofOWFicGV9VpH4CF+Q2k5JM0d5dd
dWrdVRsCQqgFjNmc4bKqnaNKYFxjEzlnoS+LfWtG9uNSSxYisFOYeMqaFHlF5SSQCkCDE4/GPnGG
dhNEympfiMwUJv3Z27yFpoJlx++PmvPKBnxrgl8sKriKdEbBeVOlzXbAim0xtSkKUjiaKT3Tb1nY
vzeV7ip4hBmn+2Xlav9d8knDFlNhwAMYZppXtQPidBntr85kJN1AMciLPNO9ZICdBsp0oIFqTiUZ
Q3+fZgczzE5twaDbnAYT0BMk3NbMVX/W1kO8dePjUEABEZAxpy7rcZJ0khQM9USq6NroDnK3b1QS
jL4UbPDT/ReXsojRdckR6SULlSx7P29jubqr18KK9qgsUSmPTwTbKM35UbkfBh63KYkLgohdsSgp
iE+LAmLg6XZecrsdPaddCcE6RWB6rhilcWG7DKMrs4STKCdWjuA7Wo2RcncwS49ZK3CXXUMlPnMJ
BMFxJezJN/8LbR0yVMQJ2Z+jXSexnarh0i/XE1W+twd/jJLXVljEESeBsolvoN5NiaEDtDFr6KDX
0f/i5GIQoA39EAQSJlSKkV7qics4VRiqulzqtjcKYE1T4q6KE3m/pe9sHG6Ktp/vVmBAVautL5qD
S5rtaP+lEUerkULXq5+4M+t3k7MFLvgDXoXOrSPkswA6/YxJRKhOIBq4aIHJiEMX3xJ+L7LA3k+L
fdCc7LQkhRCKros1s99UddM7h4NahAjcr0ldn1+kkMMQAG0rs357WzPbFLUuuGH2uSvT/52P00pk
omMOzECVA0j0adL0d0oQjxxYfJ73xa1HIWtjaw3+ttmIEutfVm8IFQZPbPuaika92xEIGOoyvYN9
X0dLOp13b9SM4PKRzVnwhrVVnTm6a3CqCpPSYgjQ3fdAWlrBRji8FtXBauqTxDscMcOCEIlPwioe
jL+gJGdpVUwNWmCzV6oO/0eAIGea+oxEvc8rDOd0B3HiEsEcjlI7iBANgSpjHS6DGWrlFqX4jsn+
8bf/vwSwYe8PBMke+kAW9wRyZe+vaPROPGKZ274dZvwLUfJsH+PBxG03kpOVwSIqw+flFPQWVaQ0
GE/HRP8UFA+0smMDWFzjYq9/1TZEIds7Kf3kHprxH+OLdaUTKtjcebUrjS0nDRV9UUSe65W7ZarM
MS4mbEFJ4YgY/2H5GU4TQF95dcMNKls9QXRvRbjH27dJiNghOGPvAjjZOBi29YSiKmqJHi76awD+
cR+sRMI4k6NKtiQAPiHuyh3vS6HlK+vGv5wJmaMMZKN8+N+7EUF0Hlfa4bVuvbNrXxVtD1jkPCCe
SSb6uD05tD+te+HHiN2+hTruZM7qrctayVuFQN8yM6spudmDjZMuSHJP2/pbVU+Ct879qiFXjBHy
kBbxjnEkQgPLyRxXknvYgEht62sRchTCotIMcXQdwU49lqs6/Ymfr48duOB81SJqnUWEnK+08JmH
ethqCKrEBXn+pm66Sv4wRTcMz47i80LPQTVW/suwaaruTRV03saY6eEXqrJErmGXaM5RnSDKsPLN
siM8RPVEdm7/3oBrRYEakwVBYNolfNJ1+P3N8N4taILpoTtnFt0Jf5ctaqXdVYG5NDafD/clMN20
3vcGqtRNJzVvMFa/OYFL2mDYgh09VeG3gztZWaRU5XV7EJ0GrlclzZNfCv4i78POE5NFoMnhig32
GlrS7wwKpyaWglBbwyky608Kgmnyg9xdD7Dy3mgyJfcOd4zmv94wzxvO3Q9jFfQ3Ae3anVB3ursG
yuMtteyIRBAc1v/PghUv8zMS/3FmalV4n3cpCa01ho4truGI80hLu6pp7sYMt09XqqhelZN4z99t
vlCx50gh1aaaOzsERmPL34mE5DdFPkut8WLNjgl/4Mm4vknCaRc7lnltVbrGLizEaJ/zyhJiFbGc
2ZDamUlB4e1d8RqJ0+Oe6kauuPI1ny5oMwn9dcWNKxhbLynz+rg6dauU2YkUfbkGIbt8Fl1eXNFp
XGgd/nij1BVda7Csod3KRfrJmkkMTxIvVIjjKuO+onWv/uH0ynkckHzFC6D919RGvo+LiM/CpAZ7
BBo5CtF+kGhBDVckvYBkc5I63koJgHyPZG6fgJaBXcAEGzp7BuZJm7N6DLuM+OmDqx5EZbV4bSQj
LoK4PnuNV5hV8w7UmS1rlBps71RJekdueWJLJw3yHP/VtVvLcukOJoPhdAYLaJNiIfz0v+L0lHXH
A3XHZaADkQEzLeu3+6n1CGUh6+aE+zPSo1Fx3QCfXuT9mycSImoyjCRK9BJ0PX6bWClrYCvPVgAw
UFTIhzACNq0bRwIZqkNLQt1s6oBKrhDWsweqKZcTQOrMbv3zFNU8wHav5ayPAiID+elo2Km9IilD
jFWvvqb2BhiOGySwbFupndnDfEEvI3dkYQAiAysiYtSg8vpHCDmyxe6ZjnyrE8zhW1HpEJge7t+I
MXPuQKnjyeOMTwDvJAYcZrb3ecQD6CHJmxDEmV/3e5oePksrs0o2Ww2dzxpEifzsecnH/3hKN5WP
4eQyd1fTMGIPVIbi3HKUwCtKyVAxQHI8xMqMNvyvuFdleN5NVbSG8h8mF0ObaJ/Dcs7bIm08Q09N
DF7ju89IU8mAMJPSQKZ6jAGL2AbPI6fqcerhQD8aJWGkT5QWuEa6GR/6HQCDpXV08UkuZXc4AaQ9
K+MiH2jmgP8dRMdkNP0GUaudQjmXp4WJKYgPi1ezE+tdVCjoZ0GfT2yQYQStA28cW5ySbRxfvL+z
of6mnDoRSjHvW/U++V4w7p87PpY4p0xytms8RhFfP1kl6QY4vd38V+CvoYaNUw8E9lnHzVygYk+O
lj0I6bN24lhiQ8xGVjwEgKJMyvPM8cJoNELBnudpQJf9lTo/puZyD65AAQgIsJSx/KiZVNh+MHAg
S83tLC1wPUHNeNOunErpvlkVE2hLLoDs4nHUyJbIuLwW/ze3rsNLcV2eMOV0NjPEwGopwWsw7mkS
y5BgOe1ahSfE5kQJYgq3/ATdCP7f0VjN59GB+jkIuHiAsaSjk4kB1dCE8i1BegHUveoVke1sY9uh
imtJkiGxhpUKKg6mv/n3fL6ljASwSGjqVzdvxut0oMwUnrbhU8D176nZw0t9Ieu2lVpmQKXi38JF
2rQFrKU+mFQ5UCxwv6uUcfYhM3kqksEmVCcfWeh+def+HV4QEj3BzYWRhsDj36ljL4nLrCURtS5W
Ko/SMsYbxrntH93X6a4t+/W7FM4RQojrWrtpfT3mKveUmbHpMfZ2vkbRb5cHYL8ZWHB2/bcoWX09
CPauVgGSTr8US0qGEVGdPZMZHPeZxU3eEmNRSVEyXGf5+T796FK+UOTt+0Zh7Pf6CyXsGcv1gFcg
Bee7E7qt7l4PBpaOX6fxzG4ozy9V8VFptH0JVdMIbinXP2Y/NuliUBw/+rguLjSFwl5RYiqVHITK
hDfxtcU1FzIn2+Hs7uVw3jN7XEpXOCFrvApihJvY/VuVK8eSGS761YIhN2+qw28upSj3OMiNPE8+
ktEZ7mkGEOTexZa+Z/D+IbKujC+AMQml8LG2Q/PLLeigqLpC13IZ0VB2vlxBqB07tJKlvcDNWAtY
cHVycYhmEK12F9gqalynBYEp1+vaflCp4uZz1ZGWYDCkCFYfI3x248SEjhYCQ1G8wOMbtAHRLZd5
+jdzu+pP0YfBcUmDz/ev7Ltps51gPF9Ql6NDN8IXYLfsmBQr0jyW/azYbaCZTocA0xJxDmELK688
l4aV73SQ10sYp/wypjDUOh9H8injga3dNzpPzEjedvnejhoG1e4bVpyjoVej7s6WCFQR05pyqqa4
dEM6kpUa9zABs14boio4JIj6QXoMGEdK+Eg0nkzTPtV2AL1FS9wSP9Rqxuua9m4TwlXCkzlBlU8y
EHevrLr+5FE7se/EkYX7b0n7ZRVzpqtBa1t84kuaTXPXb7aEyyI60Gv0kopXjja1BgF2dYsCt4Ah
9W2wVTZCuP5xNekxrMgu+AuRuVnVT5IF2mm1iYVRAWASOc03qcgXxm9wIuxVO4N2jcA+DJnCW8B1
XXcAAjTLxo8QKntauSW6FonQAfGv3Bzd7unIsv3IwDpFKo26bQNsdNnDCCZnSCaaxNYuOf5BZOZm
6TCbhYzIV3Fz7d5meLz2by/WxhO6edIl2T/FGDcgzuA7g9sN1l5OxTGtRY38wBgkdePTbKwoKQLf
rF8nRbvDd3formH+l/JpnoWhu2cmqPQ+kcRoobd1JRoIYeG2UyH4LaBPgf+USDsQCLWyltSwSJr4
75zgKlrHAZXuKzG7X6iYQd/EEd7A6j83aobYkvOUoNxcW6T/BGsYLaT0UvusX/pz2+RBB7MimHgs
4DcQjXNaYEOsammJja15ioURv505dgwdKuAcUdGwUuTdS5puSja1kuhnMGyOs9mlC/vTJ+atscUS
BXsSt2VjxQGP2/yOVhytZvy2JN5m1SM1+plpHPiMFz/u+zo5566DNG0M0n/ZoYl0bUVreH+rCP2r
Ax3epU4TsWP/MX80azvi0i68M6QatAlJzUEXCSgiYNqoxP3FwXUbA86NOM/IReokgMMTYghpas7t
RmDJXVFC0iEt95FJOlvLFG5aioDGH7DbiCchKGEeAjGd2PMourrrXTVQEeYENB+slv96zH4D8JBg
lq9/4cuBZjwTktfkABPRS7ITvZ91GH2poiubIIRbRMm6cxADl0GQX0DqpzuGq9M1QsvzCmYGtPqq
lXx0dz3IC/fSxbfipn6EMo41i0gjoVb9ZpLzbMp+sT4Ei0zGnm8pALSRuARnlgy8za8GJjmtuZpg
2Hx7wh0vi9x7YGimtS7VAcsQxwoMcr9cZCBTTLPOcX0YjDJ2VYgbEMP6IMWkPhoWBawTkuXF5JSJ
BifVLVGkR8d700gOS74pYsVKfwbe4bcLKdACQ21JJXb3o309PP8NE2PLxrw7T++NxWm29ZP+X9qv
un+n+gIt7zxkebbiiVY3PrVNAXgNj35l50BkVcRhMDgRusPA7RawHt7JeGDljwuqvQm42KwotCko
z4kovHJ2bdzlL+7/bBHiJMrxQxU6mimy265+/1Jlwn/Gm0jeMOyEF4elQLkrp2WMKpTgy6Q5R192
HQL7cFb1bRgdlPbODale4e8SCmTIPQbq5Vf9khitbKFlfCohTNXxX3JVb0GT1AufeMxD/E66knPd
kooeE77A4mU7OxPEFAq5JMGKObLCSr1BBQ6zcs3gPMt1JT+lu1blLUuJzUVTeVo3AuYP/f8iazsV
AFl5+yAeLqTlSxB3AsSgqrqV5m4jhx5N4xqD+TMHO3A+jF7sH3lrX6xla1GmLgRCtoaB0MLWRTHP
7SL3vDRoDImTtwFHSvhz+xwt7UmGyv49Q4MNjABevWT5V1VMp04Al4TBg2mlQ+K/CxRF9l8qI38S
FgsYmU64Ozq5l6CaQzuhAL7KnPrMqcUa0GxvbohaVwcRubh0FHRH5mreVcRQkxDlMbqrA6oDzex+
XPErQSIB2V9Fw6cXRVOKmzN851uQE2pZRULjXSyH3NH2fEoOI07T9fjnssbE4AyjWUySf21pp2QD
Ui5PoYejK5kMpQDCdTX/8AuNF3XXjSDh0VJwue+uEDIqYeK1cRqqLSC+J1vfcesC7GNi4LD7QuTz
vkNoyAG1p6IjgKdA9I3UpRBfByG1DqfnaLWsJS93CEiLMfYsCzuOZw9YCwcEKs9uClsHzf0ZA/Ne
pWkI+10x/TsjZKqS0CACWseuMKo86GEhtB/ArMyq+hQ8Fu83cJhrYblxN7ZF6+6cQLCAkRWruxfV
zwVgBLLv0G6KfYhIyVkb0KzcL1mupCDDJmclLIZCv+10a9d0zPjrUyMkRK5ylttVL8FcY8cDV1wj
eYcCMCFGSPIxGdI7KkCFfZ3bSTTxd+uxqktg8p+1x8NLueEuoQhXsh+KefWei/RR+cHNLYT24cVX
ZHw0tVfpqrp6s+KY4i0Pt2eS+KJDrk9ueJ0H10ZhDgo0cJ0MF9us2s7lUoxkl+udUktTo60h94Uu
B6GuIRQo0m4gGW1GFTPrfu/ur/89Ist7tKsjw5/b7MXc9Kdx0hJQsIhQxXZvyNfqq/IU1AftpVpj
5q5nuqa4C3VbXXj2WRJV0aoa7chnsncZeRdujcNjPZJ6KPKc68EmFqqSdOVfPH5f0zqSOSQPEbZA
OJiVoQzCAXCyeP8wgxOMGMKs36EebYpP5LL6TAhn1mnkYUTgsyZ4XhTlHEChW+Q2u943pPmSCvve
1rNOLcu6kaGqPZzgvNEb9MFuTfKWh1nTaZdLgreIS7WvJMofXRQ+KHQ0XEAG+Ohw/BvMRyHn6lS4
auLlgK2myQpwNV3r4yzrgyoDcyr1Hsj689A5J9tfDJuFzrfZKaD4ARoMiwOr1pjB8gKx5BY7uvIR
MSOORN+T6C5RFf8wJAaAMwyB92kWSKTnDIzyGkVe1DC0co3tsshRbkvmMqm0YNHDyZnWP7PvQABn
D9lHk5XPlXjJ6Mv/K/j00Gsx1BpmM/xIhHy5smrZBbp9dhmsMTyq9kQjMLfAcRF7O9d0Wu0plWiz
4Z1a/MRyaVSl6w7vkFO5UYSD25C5a5pFn06AlINP5XbQB2Wp/Mjm7aMp4FnyVPtS+LFvk8qT8Lta
Qq87Tz8dwTDAmlxcXR1c5Phlh4p6vIbB5vI91g5PQMScQxNtcVVPbj3uzV8nbF4A/6gUhcprkr5R
d+eKTLI1+ie66KCoCCak0t/wxZqHFdMUp/2j1gOi110azStETFEwGJPD+LAF5uD3buRBNmQokcdZ
YN2Cy02OIPOGZtzv7VlKdClUBX/g2oWO1mfCRkTaPD0HM09gGuQJ7sfxePGsPRPToc57OW/4FwRj
62BnJndVdwvETgrncJ46PneBsrLV0+BXFxiLzglmGrGQG3BKF4c2N5R8Hei3gAenVwJF9lC2tUJD
hiCqxTPLezUM/PAC2umKtg1irmecwW2N5SrH5dwJhaXQvM1JCWhm6jCoZfo+z9Pdq+Iyj0uboBY9
iDm7fNweTBuARRL8cClglS/WY+FmQbBl3PD/4chYa4jbN0a/t78QCBn9abdhxMxRwC4JsRficbK7
q27MN24mcElo2V++YylRZN8lBSep3bYAFS/keoanZ8Brk1PSSZIDtF++MxYWaa52zfmkCHF/fLU+
eRVaM5XmZGIJzR2o1BOeL7L/jIxrco+dGMLTb/4KDRpaf6mQ2sA9SY9TEWT0uPIomPN2He0Uhvl6
ojMUyt584Bk2ejOyg6iW/6ImHIgA8WQnapcOi1I90PRUGg87OTQtHft5P78NYVIeXtckVFTf4MSb
Bz6Sj6e/VCT9508AE2y3tVpDw5bTBX48GTD1iuWBaW49BJ1BoYGZeg3MOd2XIdVOBi9W0AzuqY4n
FcbUtdjTjf1WLqnA0t0pxA/9XVPKfPIWwA54yZiLP1LX2Du82TWt2k0Qx0N27/fkVi6sMC4tcCJr
hpYQfICYFJ/aG2vA3RMUZ649WxhBH4XZnlhVCDG8PufA7EUwfKoWPwHEhatkWxfB6bxS9GlJSM/K
OZGNQP+cZcjKgRCCVVRmQcMFygnBJaVv24lVbqTRsIaJ2m3r0gs861o3ugrauNA0vVPu4p+a8QPi
sNdoCRiFLtxVFc82qC69lzAREJvD2G+7yPgn6K3ifKmo9eQoAqjZ5SG4A6u1ljNhAXzoIQI/lR8t
U4pI/e5mVxp/wxxQZHz7buj/k7ZgWk7ovkTbOy4wk/uu3+VCijtb4lzgRQq5qTEeYeyR+Gc3IdVx
wBdfvIW5A/cb2XxfmoDp3xfT5EB/okc0qc7nhXBl3h569tViB+XiYnrG3W6x1EnPrdKrEv5MGro+
NFpvKoXeF7MCm1CQPZ4M5snr4OpFP8W6w/YK+Fk77q+VCne64VsRF7xuyDJALTClBQsC9n5HprE6
oBoWPShUi4Ous4BU/WIK2kYBMnty3k3JhnR+GcrwX7K+u1xtFOO3EHXzYbRml+qWMDXmCJG43J2/
Vsw7HzKYBU6kpmtyQV4hKAJ3SWk6Z1Smz/geFbJCUZEM0zVSiAeoP1nfLfQ67nEc5bxp6cjHNlX4
EJ2jtQrz33SxZel/LIeEtsO/b8Cop1XehcJw3bRv/RyUoNahX7BWwWkvOb0ppPVOb0B1YcbzvCqu
d04iBfbj/JUFg+it9QxpoNjpJOJY2FgGVMQq1Lte1tJa6C8ba/YT/exa1wHMO6Z7H5odbtJx6j2q
NGSrzPMlK3D+wBIKw5R+rUJRIO9ILU6x53ja9a8NV4gaIJlGKUNXaXinIMssrjaihx0f4H2ZfYmi
ghUb6A7yNpkqLuJmAOuuAwF99IpGvI9k4EGiNG/aJiz4BNUNqPRzlcyfEoquui7nkT049sFpsb4H
zhLCfg1Qp3oNJMmvgpsehCMeudB/OcJRUYuRF2kGtgm+7sbmZjGdQdpoH8CrW8g1GhOcw512pAOm
7q9pmdG2ttK2N1CeA7X2eR+boaOHtpyKG29XCgvulAP03BSplr+K1SyV1lMdF1duIAAf2/5LKcVu
8dYtAUxHu1C4SV2blbcVPhmW6Gj/rs6N+ORRadoI+kTe5MqWQrRP+/i2sUrHxpYXgmJBWwe3MAW9
IxkAzdhiTa4sQLAuEah80Q29dA7FQHo3QtkrVqJmpLLu9xC2UxXoR4FMDj/wjpyu7clcAMvtArJc
QG/TVxPfpfWWJmU5KxAscs4F7hUUYxQ3Ms7+dnawNXwJYZtuENYLfa9nrs6jcy+Hv1GqMs0cBRn1
fS4CsciTzvHZfopzTi7blVKQiYl5t/Z+LOzrbT6QJXMdwF2PloUCWzn4ywmZlvq8Fm8O3ZYr626W
3plEzwu+X213t/ZClvSb5ugwPtY6mGZPNkJkQeZG907E0PMSNK2OEyofQQsUzgHAf3x3W7HSFksP
7LK4EK/S4/gZWfMRbh2UOvrNesf+6Ej+euh1uu5Ypy1hS9Y7gZ0Xq/jcTUJ10Ce6K2uOmRdX51sj
LavoYsg6p4g6jFXuIrWXWW6XAp5xxSMeRuZJKRyWruIparU5yAUvn6PiM6yOceB1cxc10ypD7s46
DTljOgVGjjxtR0NyrNRUMlBH0X/+iBmR69/5Vwi8FCx7AQi6lDvLosxiMz4NyDFJgatEP5GbbgUh
/O+rOgTGv4RAw+8RHuJ1axhGk3fW1djChv4BfQ0XlKULk+i0AUrU0fpul68kd3hhgkcvsK5xi4OM
hsze7/rrncHv+blsmOQ2GRqgnVpQmK5wwooLAfxWiEsOxP+kvphWLfKFoD+J7U2tOliuPJUMdfXN
rsAAd1+WZ/0AkaggOZoT2LcftnIstL07rfryGh4f1FK5DEx8zsDLAmYLktalfsK+DKnfGsu6J4a6
rui2jIqhOcWeRyY+bWFu6VpwyGWLnq3Sgf4Y/niOelcXfW/2dUKoa003wUhygwuzgiyICUcWePPb
FWmQEb90EDTdGGkpkqMh8E5t0WG6Dz45Kxv674nBJzU/+pb3fc5DGA3g6MTeOpTqjRdI2O6mMOym
pRhmzkLHIewlu0IZtbGNAg/r9LRFpJo+CZR+iSd/fUXz1YO/OHuqmtB08wO5O1gapnN0pUJIsFcl
bJkgAfSOGaKS28SoKYpCr3Rn31H/offPzzghdlhwjF3z2LSn+g3+E6212jpIftfy+KJ/d0tYqiHZ
2iaPz4snOY948Zgvg327GKQsn0W7n7xC5h2MV372GfWOvg8HeDnqqspjHDEaRTQudIrlJ9lPPFR+
hEXqdr4b/VVRf9u/yQgALfD5+iqpcuSWdft98rlCcJCAfE9x/1dVmw8BGUsSVhXf8Nm0dazuAvQQ
3SWY6qWkDzA4woJ/CCVWXhK9hDcERuQEaP+/hLGFFECU/WGFAf08iXEaAX3ZQ9S/tCX8pg/T9K3g
QonjhYHr4sGtmZWqY1rGgfDEBdnqcEp+SwRBYSJCJ/0DglRp+KOkhH/LBy+JidVrIX+jGuGTsg6D
2jMEpcZtOPCj4Syi64PH8h7YsiZAlDpolOh4dUva02c3gux487Tzbj4KbsMd9yPnqWeCHSVNYlit
HeRyIEtcHzCgKishGH8KzbQ7yDIXdUxcD02A2U4f3uAYF9CHtO7tpa/aMqKFlGHqnDVYqXC50oEU
/RLb9rPwOCZ7BFsCyBhnh/JxwehRiTAx8caKTRcliAfiBTa24vM9rA5d+bCvYc10llf1MaB1zPcC
qmlNnajOnZZ19Aqhx2uElVnS4YVcLl4f245TKXtNV/vnan0KKskErE4NNsBruFzr/WwKgHlCbR1P
FsfUY5tlGomm/wUcDdf4fZZsfMXe78WzYnicBbB7lLEAgkl3o8+4Kic6Pmd/A+bYLcMMOD5o0hVr
ThmdKUcMiW2No7wngDRAvLfL4P1IUUgFEOJAs9x59QsV4CfOy4Q0Ga++Zg/K56HhTK21Pwrb9piK
pqFNhmxCkfoHg0nslWX5M65TiEY3Z0Ac3SZ8qFEv/rGoAV6FHUdqk5wG0S+75DdABzaEes8zIyCB
xPvdc8xD8zTVOkOrIcdcFzvtwEFIgFTZuo3RdbFlEviOkPAv/PYe6VX6JBGFH2Z+8saBMWY6fRQv
Zgp4dlMDONEU5xT6soL7pZ3mpbA4ajKQZrEheXSB9IkJHCXXXCs/fYzvkWvH0cX5yWjCB4ES8C2W
dWge4PTRyBNjtNuH2NATnFcJ+NcWo/WjP+Ze+WVxxb4vmGf7iHl4rLalwUidaJsgs4kM79C9mpfr
7deaaaSu5zE2iqpFN9lDBS40Bc/bCuXnL0Cpp8lPEt64OsWWxhG95jYketL6OHFL5oYyvmHPkaeI
NGNdEMnIB4kKNtz/bI/KRjeqby6ZtEX4/sNEs61UC3clY8jbFRXoNW6h8jj9n5cpSsxyDi4z5rj5
b1sOkqJY2iDFtiJ6PCi90mFyFJX3XVZF0rqUnRBnYYXJ80xv+PPDWgR/NRNxGKl4axUxp/PHlSDz
LcS1oG1+a0AeGBvt4EnEEn266vtUlsU8WGsBMrOsyQsDORrH2d2NxnPEBjsNZ6hXmHFfzjEJeTbE
GfX9FBywyNoR84P96uES7krgBEi2iAx4EFekIPFoZ+8NI9IUNFrUz8KAt4hkoExqtw+eLIdaU0Et
XuxyaTEknmG4Y0R0D/ZIqgkX31aPEA2aQ+NSI14Zn42IlwIeCI/buwizT6cVvHBJtkmeshs0KJCQ
MiS6SzARMgelVcX6ETHZ1v5Is28Bdl9CnKi+ZvMZ4gRy9mJ1FUpYeBdwHehAS8z7d539kWl/zDIz
+VjBajdn/Uq0uwYPCbG+XQSelBVr0sL6lipi8vfbYw1zjBfmoh+aVAYe0j/q+ETdSGjh1CQLAULV
HFGPiLz+g2QYoKuonLDg4BYUNDkkh2LCJQ2F6pPL3IfyRsCZz3fa0RjslyPrkWMzy/rvNGGuWZlH
Uj8h6vLtHLpMSNroi8MwBxWDv5ft/XafUFfeI9yeDhgQsU9Y9EGzBD5GC4oU9Xbf+Qz+LHbYEODA
DNkri/5IfvIcs07QyXnZOf4z0QpvO9m50/rpBOOC4R4TCxVMUlO5g5eHrt4zA7P8MmNX4hAAbnbv
kUykYSbvsTuWa1/ymb6/ZlaMkMwOqw3eZXplmZAS9t6WYZ37sKjbpMvQctm/Umsa1gQdtUN/Nlrl
FpGJM33gtAiuHM9Zt1/drxEPjPNuQ5aVCtbqEeL6dSNGEX884CGdY6IaMmS+5VJmeZf+OIndD8Bv
y+QoZGdhgllckDx1z8yDitshaXCcABQpSdTFSXEGsNDfkfZpcI53iMhbkkvhoI4mSNO30oSL3rF0
mN1yXfB/S/2Xgh5yOcNOqKbMb7mLIyj+xuwxHtR9JZFn37/5n/32eJ37FVfufs0A7sygE6wSMKWP
arXbDmQHbM3iDngFdctpUC71VroQ+yf5fVqYnc0MK3Ay8WTH7El82iH6A2ky4X2PrZDAuAtZ6E3n
LWa24D5nSPyD8ww7EfiEqQ9cDO1U09ptW6tm339TAk/bui15Vgi/MCf9zPB44rRiJlWfhwAHUv22
WScCdJwWlLXqwMZuGAlJZD67xlT6rnokr4uWvZ2AXrcrr04BUfjH5fpwhoEpVqcw/1vuIfEMGVxA
3AnON1DNw2KVoHWxlQeko7je2y36US52bxGfU9Tf02c3QQrOemS/D6nMeLV8SG8JGOFp/edxW7V1
jiXrbSnhndfJXjggYuNzNqHmkQojO0kml/6H+bh547yRlu2CNtlHu9a6Ld8ftYdkVU3ulZGZhGIl
NWM7Z9EaL4nZXyk3DDhlTvHVwyCyGDoTiqxoVZbWFX+CXbAbQvTkkyhQfFp4fPaZyao4VfQAc8eO
jnv4nedfel1OVjvS5PCRZKowwVxfsqB3WZyImY6sA9X8Yh20I5KSWrB1h4OKVr6Gvs6m4VHdxG2A
Wp5jAaIcbYCoCHOOPcTprLh2rJnXARQ1G1f8bDR5f6HeCAXigbbykxhyrGnf7iqTrtU5h/SSxPe/
RiiqAWevAQysyY/p3gIKw/EnI1WZSNIXoVrGFgD3tzokD7TGqPCHalGumWxAS+JICMtdCXhJM9lT
zAbFugcBkgiaccG0TSS1keF6HlVTcsFC3IeZJs5//t2NbyUgSlyrppi7WYB8tI50MPMvKTaBFeMg
xcsDCTgE5diFZHz6F42TzUh8HiP88sVqPQsPxbCa3UqzY2Tk6wmWfOUKGO0405kQ0J6A6uIUDkhk
v0AQG+FgaKc1ti+tBB5fCYHDILvHf6kNr9B0fg3qv+LJtQCa19BW7qLank4KiMWmnSiYYPx7EU7e
RqbHyW9du1VnkOoMUU75RWPz1KnFY4OMCmpAkmzcpET7Lvw77dbp+gJsau4iAUVa8PFF8L/1BgdW
wYPiNvpypFlfFJ+zEdMfeAReyZcgGfm/JKwb9/G3v7llOi9I3+kGAZQhr2/QLHqjHnFQU882rxZf
1JXxz3979HfsstaeE6SgFHtA981lj4Ug5AxGkP2e8Rl1rPSkhTkz43d41aADcMrnUVQMviSMVRwh
gP89V7368Y3wPqZI9bQnlgnvGnGlctp5aeDRAiqy3NNP5zwRKnTcMjJndVt8nq+N0CyIQ5czukSJ
75r4LXIUgw57Xug5LvqBcJfFGo8XmSEcrhM8vltYa19oLwFPTjWhMB4J8BKVC8RnJA6IGukQEvlM
qZsOAEw7RSxBg1xW7b/LDxPK0c0pezaq8lIN/p+b2eX3MiBDHcG/5g5Mx0IfRo38VhtCF7a8NhO8
q7hn24Mi4RQiItoCWg0HDWNjOUuciMWSPW1lVMFFn92aAbnYs8xejj9YSrWHwdTPGVmFa9qN5pyO
0Hs76/nU9lZekhemnMdm+661WI2Wvk1y08juU00oQAYl+Cg215ikvJ4o2A4C5VxhBH3sqbeHiGRk
re4teAQpEfvDve1aHQjtJWFS3h9pRbBDOKC8TU6APeQ9ueW2csQ8tgm1BKSVaqNwFeMklhimY5fB
Pxmzy36axK5Adg1vTHHNg5+HILAGmjKw2Jq8r15zxkTLmn/yXMwJSpgYIp0cmWtPvgppfpJqmQNV
kkyXpzMp8Byj5W0YRXa43lwp3XJymOTpkZpEVwfhFOR5UFBRiYvcfq1dUn6+Q5KEfxBmmUWEob1e
VahHnlEAlpfZUp773aMDV+MO4FMshpzFZBOcRoAepUmkLMQ3YxrcdjYOpJc+sdBEMJm/UQX9pTxV
K2J8EfKDxGt+5hQ50nImajIRuG8x0N8m7MAWDc7ZA9/HyfsyuFecCM1wMj2C8oqzMbX8/y8guRbn
SinkdSA2OXobc4yxMku56SU1yBg2t5RSWcLgHoS54egmoIWJd2/C9yeITxnolKycE2e8kpHJLf+O
Fm6iLtkSfRIYKI8tj0R3NOJV+12WmN16fVLs16Bo6pN3VTbsVCOJpXc/CVycWGNf0EiVsl64O9rs
8M2gc12U6TDRjbSFeHLQK4yC8R4DfPmZgw9KV8a+oIngQWj1toOxnMxeOe0WCJhB0fHgQWYwanUj
ALDskPDeZbY0QKVDNDqPwqlBjpYewDjwaq0CBiTO868eNkj0N7O6gH8qeO0Xlrz0wRgVN4fSmiQ3
TnR+TQtdIV0+szTpMTDyJ47BvNQ1Ta/WJCBjMU+x40X+iJjJIV4IhQp8lE/tmz1z53bbj2wnulPa
lGaTtrvIHdlcrU45t/pAElCelxF7zA1t0V+oDTnOB8xWS61NPW2XUm6NQ1Fbl44GbTtqf3NMtbP1
+vSHJADV9DLedMlY2A0BTFuZGeuF3mFjMY6xQhortkQAxf82OFByZ2/XUfJmoUKvBv1yNqJjkMng
jJ+SL8yowT8r1/PoAAThyC0S7FD89psVzxVtmsRu609Bh+XCnzY3cwDxwXaOgjnRuj7s2zM5cArg
nS6mXZt34w5S7cqF1y0U1oKnJKEXJoFaSAsYW2SBfTN3yDCFqdLX1sHQMwoJqwKTn6zsYUZ+cqgs
ARiRup35ZFy3TD0cZrm1H8xKkcC/wFpAX0pulDA8iMMWJWNkcJOfmBK2AvjH4E7hVgQdZOdDFDUF
xHY3fEwHn8j3wnZkg1f8FSw5SM/G9RnKUr+uTcRFCGW4bfjIn4wXTQMDwewC193vVJ3F53d6H2Yl
yCEQMfXB+YwegWjy1Mw9D1WDMKPF8aqwX7DbcvCJRPhWkyNnLSC61BrKgkgo/yydiL0kZDmXuCr7
Vym2iOu0JbcUct4B7SC4pXgtkzJaCpMbPfHFkfYsr1i/gmfiwBwB9QF3WJPmU93oyZrevGgTmQVi
t+NkAiLSHw7Y1ZGeNrr2SF9oiqWpdZjWlC3FMNmaC4FtRZDBytA71wYUV9MU/a/M2Y6U/mNXT00g
QynsimL29IevYYWwIDUTKC5MbpZyqu3cVe+iBVTDOTNHwSh0O/wPngc+DJoE3tajK9p4UvF8w+0B
qB+yYyjHYtF0+MAa7megw3fhnWtng+fPdBW6Jj1aA1rqzoxDs2ic88cmx2fiM7WfLumII0JbUiuj
BXKkGDXHvUVYwfCw49JHw7cIBBxHbYi749keZW+7rcHFPXY+Q1xnYcw6203OXTJXxOFaKugUrckE
P74oddnB42IQDEx+T3npza3nohKDTPc3sF6cn1AuY+xJ+Vk6VOPHte/7GeKb4q8/AL1daoE2Z5PJ
sBS7g7pmEISYhflRHJ71P/AZesxLMg4w/9LNGbwkedfSTiCMBKH9FHggYCw1LwbnYr4V8v+GdNHp
mYu3VZ9BEgX4rspUqcguK2j/XdpOghF2MEScpMi95MnVa3ftyA/CUBO/Y7GvGTf8VFnv94n/Rme8
ZhmGkbX1QCp+//qYWUThKcW2lkTGZxGRO0rJLUhMlrQT1HkyGV+hEMXOxsJju3HN6naz5LgNWBmZ
3hZwzFZgnovGFILDm0oNQvcEYr+peuTObBDbH6iHlae3aYRCUCycGWUJ6V5a6xHDrXq2iBqW0EWa
dkQ+Zd6hoss87v4nv3Cz/MdwHmPOf2Wxv4MdZIfglg8PBKMFJG1B3ew8L+P7ZJcsjH6YAYgOMjzr
O1grReoAmQ2aOKy9EvtYX+4ilGlJ308LvfGZNUjssYtX9+mFIosP2Q+jqNrdbugejv8E5sjRI23V
kDzdpdyqkMdrJUYsnJOkttCB/ZgEdQ/3MGM+TRl7IPrNsT0aR2KNkKFr1nE9FbPGmiNFXHkGdcmZ
Xxbfz643fQszQanWfFWPz495NyYYYUs1lZ6+XbG9rhB7cNtRMv5R2OiEvhRlvWEwD4PIS+2Vaknk
UKOb7SPYAz3CdEcwQimF4DJN3bf6h+Zn6hYj0/ZUlDCjeyUIWHms05yu2LlQhYidAkq0DPzXOPjC
W7N+LWC66Xb6DC5AH2YR/yTpRa33dL0BfLnEAKmwYEbCXJM2dQ5tBKE12+9UhzeObyAkPG6OUIGv
bBoZYCXAFMkvAPADoQwnIkm59u2MgeJAtZUBUt/karAYMMC+V77JMGSX+brAJXqYdoXXBW9TaoJ+
foX81yw2PUirN/LQ+3hJUyNAJQYmIPEMfJWkB5A8kNaQm0YxNAYVce1fJdh+xdaPwtrVJaM4kfET
D4eHOXu14YUUT5L9l8WjWY+6lItE7/XZhzVqcmbUD6149rSC+drXsThVFPCy+BtCSG+v81fM4HW7
tBqGst+K3h3vwu+CjVog0wT1dlk8NP7tqnAmo5xfBInjqDR/HlVkprkCyENZpu9euFG3JG1o1F/8
m6jnKNNgHK1PPEm4sX5o56+Qu/wz37LSWkhS2AbrdU6K4Mo6FLJ7qSw3rEXPmBLLUHFqiSCLYRf5
1IpNybomXg0RuvcwVLgCtO7/7a+00tUOuaMsV4zAtn+uHahGE8R+eriUHnxgYck2+OCPz2B/zK4G
szwf1IzN59VgAKyCtniANy5QY7C9gyGr0FPaeuCKK28Obxs8Oj+c7KMVAYQZ8tuPgbJchEpz0gnr
tmGP6NIfY8dlWRhuwa0VSjxRFBr3K/dSKai25RBCMU8TrrBq2Ro69bYJnc8vbILdSU6UOYlDoosz
tONQbHpomLyV/oF9EgtPdwMtkzBGiJDzEHtVQflcjB+1Cpt1rTcuEQMkaNdOuvzk1OS+h8OlK12x
mFcBTvA1o/GkWNoNJ1SlBTgl0pWJqrMnQPPXZmpF8Vu+YOxGNrkU41nS+qy18J78PVd9Iz8MmI5+
EsO2ID5NSRZThLEiSmG1lGUG8a0uee1L5zT6cD2boex9jZyEFwm27qgncLkdq92QySqHnLuptc+f
ARNFAVEB1wZH5X4SkpfNVZt7BJJjvcWhKui+bezA5Ag5goY+8wNo2MPnO99s1Og/3jVTykelWSJH
5uduy0wpgA3Paf/M412uro97AWvis5b/vicpv4gSIIEeHjBJslr8buWzvbXY0kK4+YEzIJVpoVH1
EluEh7iBybRziK0g2iM+qTfcHbCSWnVlp53v8Uf67yAAtxOf8z+CAusrYjd+Kd2lbhyHtrYS1fsm
7cKcwz26APthbPbti/lSWnSnwdiEhDBE5pZ4gho3MI8C8UMBbg3UBFAQ81FFU1SuqwZR44wxaA7B
4Oq3JBdTN6DLNdbcOZA28YowYhJNr9bLIFOPaQ6bueG7SbYuS3IrdDFol4XN7C4tCeY4B8K+y5z5
QY6EO09Utj6NEcc+rzSd6uE5SfJCx8pcLI+clxJJm2KRfi3nm6qIt/qYj1DxXFoghVIkEKm3fcyN
/eA8rrUoCDmeLKOC0JW2ZpzWzuLzZhYtS/VAHHoRve2smEDNjwqvKPZQXkDgxxlIjbAAyqpe4Kmo
X1EuouHrhW7rxX87DN2SpLE2LElbk510WaGN+w8C3cjboDcIr0EKkUf9a2S2S5/LCLFWMg3QA1SG
dBXHVccPUo3zzOWS948p7nlQihIDyjN5AyFS2bL235fJnPRwUPSCemnatT758lRWuEh9KXRxokGC
uqz3LSzNi9YPkfpIhkktx1VUs3aRwdSRqHAOjp4PyQD/sqRWRH/1NC2yNWm9/AR8wyiK8nUmA5SA
mSUHSJd56eHD1JFIOShT9/Z82MmNjZddMdDfRJDrlhgRcuu7ju/SY634RrEksPyKrp72CduDwlxg
6BV2AXBDXpGrtr5OoItiM5UYQdhUIxWqHPqoJvSS1pqRXA5AjIxpPs9BPIV8yRgB+3eBWebb2Rz3
mdljwhR74FBgayNcHgTaIcqqD+mPyJ1+1SPCSObJrQfVGEKHoDrYaT1hd3UqCvjSDo3Xz9SXLCFo
NTSWzwNyLSXz/ThYmSjsAiftzxy/0SeBg8Hl6AO47nMYv9n/fWPhZb17ukp9J5duGSFqfC1XmD10
A7ME8eIYOeqXFNx+pnTTF7XIhhrLuFHdhGkadNhsDi9wYwI0UYJT+SgBWni5bk6HlS4vGJm+wsK9
Vm0qtmqccH+xdv19mLaBZTppkTtY8HHsLcu2vLneQS2rpRdA33SnKUIYIRWIyFjgP8XAyY3Ho4Zg
JK9i1qCpzoLANpGdZ88KaEhDlRMnozcU0EVF9MxEM4A/gieaqBCwv5p9MOGOF1+hqQHezxc4dfVd
OSGHCLp1Yudtz+2Vjx0YqSB5mGOIdZbqz/kwD+VgsHdsCk+E6Maf4pVFtmSt1FkeqJ8Am8jJAjP/
kaD/Bxu3/Kh640/CWf3L/MroUthIuFLIaWswcvM+eynklWcjArdLDCv6uFDfckS6URN3VneL7VGg
sqEiQTfaktUBj+b9GtJOHHXo0U4AjFVXrvdIZ1XayEMGHm8JYwXGju5h7a9BEv5hJTNm0zqEQrkt
0k5lTN+rE7FetEGtv4gkAlI5WsH4prPlZkk92nAkXwXDVddXjMOOcDcfhkdj5jm90vJxwWc80zw6
FndstHaE7KuVG89gu1AEJBKA0KE7t3DejC371ZOw6CyntbJkvYnhKJwKBfG1uwUgDbA5P+ahVr9p
CcBK8QDzHeCoCckf1UiothOL4sEFrA/hVqV57N2GrdzrjaeiMOZ+KKw3J6wVnK04eeAHuJV1hzdf
+vuQs+taMcgmFdsBaqSuhhP0BtyNktpQDYjRmjLrxNHG/4kjkYFRwFFMm5brHP8nIh1jcCfb4TVa
Oj5+0sSghLW9A9zka/5dvw3SrLKjw9GCfWTxVLPE6AcV0QhKbFTNtPXVojHsCxjJlg7eyqj4UbWR
pLCjdNSXbd/XASDbMuaifVWhx7BTyvZnWoFxN3A8BySXrZ4hK/l+6m93Q9dTvxI6dhe2aBSvfr/n
kQ5uktCB/3BySEg5wS8T5nfn9A6Ucl+Ddi2HOgqJ7PGHXtOGTu8PfM0dhLho+2WDquW8q18yX/qJ
KOMWbv6eFnAHK9SgGzrqpNyNfO8l5DlOkExpavXRsqC9zJqKaYnd8sP09qBZgC/sp3q/TtTcT3TF
1JVQVW4ULwWfX3FiD8Ya4NS+XxAdNXPl/H1AeaAdjKMvSu3ex/ocS81KR0LjOC3TqLgvQ+KCVj