176_2239_12_14�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_12_14"uC^6  �@"��l7     "V�6  @@"uC^6  �@" V�7   �@"V�6  @@"         "         �
RAM_reg_2176_2239_15_17�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_15_17"L8^6  �@"��y7     "ńC6  @@"L8^6  �@" V�7   �@"ńC6  @@"         "         �
RAM_reg_2176_2239_18_20�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_18_20"L8^6  �@"�#6t7     "�"06  @@"L8^6  �@" V�7   �@"�"06  @@"         "         �
RAM_reg_2176_2239_21_23�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_21_23"L^6  �@"�i"t7     "B�/6  @@"L^6  �@" V�7   �@"B�/6  @@"         "         �
RAM_reg_2176_2239_24_26�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_24_26"L8^6  �@"�;X`7     "�V�5  @@"L8^6  �@" V�7   �@"�V�5  @@"         "         �
RAM_reg_2176_2239_27_29�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_27_29"L8^6  �@"��i7     "�~6  @@"L8^6  �@" V�7   �@"�~6  @@"         "         �
RAM_reg_2176_2239_30_31�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_30_31"�@6  �@"�DCW7     "O6   @"�@6  �@" V�7   �@"O6   @"         "         �
RAM_reg_2176_2239_3_5�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_3_5"eR6  �@"�F�Z7     "���5  @@"eR6  �@" V�7   �@"���5  @@"         "         �
RAM_reg_2176_2239_6_8�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_6_8"L8^6  �@"�)tt7     " 16  @@"L8^6  �@" V�7   �@" 16  @@"         "         �
RAM_reg_2176_2239_9_11�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2176_2239_9_11"L8^6  �@"��q7     "�y%6  @@"L8^6  �@" V�7   �@"�y%6  @@"         "         �
RAM_reg_2240_2303_0_2�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_0_2"��K6  �@"�Ek7     "��6  @@"��K6  �@" V�7   �@"��6  @@"         "         �
RAM_reg_2240_2303_12_14�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_12_14"�]6  �@"��Ko7     "��6  @@"�]6  �@" V�7   �@"��6  @@"         "         �
RAM_reg_2240_2303_15_17�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_15_17"��]6  �@"���^7     "�)�5  @@"��]6  �@" V�7   �@"�)�5  @@"         "         �
RAM_reg_2240_2303_18_20�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_18_20"��]6  �@"��'q7     "�C$6  @@"��]6  �@" V�7   �@"�C$6  @@"         "         �
RAM_reg_2240_2303_21_23�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_21_23"��]6  �@"�|�j7     "�'
6  @@"��]6  �@" V�7   �@"�'
6  @@"         "         �
RAM_reg_2240_2303_24_26�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_24_26"��]6  �@"�2s7     "}�+6  @@"��]6  �@" V�7   �@"}�+6  @@"         "         �
RAM_reg_2240_2303_27_29�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_27_29"��]6  �@"�T�d7     "��5  @@"��]6  �@" V�7   �@"��5  @@"         "         �
RAM_reg_2240_2303_30_31�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_30_31"�6  �@"��xJ7     "G¦5   @"�6  �@" V�7   �@"G¦5   @"         "         �
RAM_reg_2240_2303_3_5�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_3_5"�Q6  �@"���V7     "G�5  @@"�Q6  �@" V�7   �@"G�5  @@"         "         �
RAM_reg_2240_2303_6_8�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_6_8"��]6  �@"�w�u7     "��66  @@"��]6  �@" V�7   �@"��66  @@"         "         �
RAM_reg_2240_2303_9_11�i_pcileech_com/i_fifo_32_32_clk2_comtx/U0/inst_fifo_gen/gconvfifo.rf/grf.rf/gntv_or_sync_fifo.mem/gdm.dm_gen.dm/RAM_reg_2240_2303_9_11"��]6  �@"��^l7     "�6  @@"��]6  �@" V�7   �@"�6  @@"         "         �
RAM_reg_2304_2367_0_2�